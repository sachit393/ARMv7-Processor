library IEEE;
use IEEE.std_logic_1164.all;
USE ieee.numeric_std.ALL;





entity shift1 is
port(
	data_in : in std_logic_vector(31 downto 0);
	select0 : in std_logic;
	carry_in : in std_logic;
	shift_type: in std_logic_vector(1 downto 0);
	carry_out : out std_logic;
	data_out : out std_logic_vector(31 downto 0)
);

end entity;



architecture arch of shift1 is
begin
process(data_in, shift_type, carry_in, select0)
begin
	if select0 = '1' then
	carry_out <= data_in(0);

			if shift_type = "00" or shift_type = "01" then
				data_out <= '0'&data_in(31 downto 1);
			elsif shift_type = "10" then
				if data_in(31) = '1' then
					data_out <='1'&data_in(31 downto 1);

				else data_out <= '0'&data_in(31 downto 1);
				end if;
			else
					data_out <= data_in(0)&data_in(31 downto 1);
			end if;
	else carry_out<= carry_in;
			data_out<= data_in;
	end if;
end process;




end arch;
